library IEEE;
use IEEE.STD_LOGIC_1164.all;

package control_fsm_p is

	type CU_step_t is (
		CU_fetch0a_st,
		CU_fetch0b_st,
		CU_fetch1a_st,
		CU_fetch1b_st,
		CU_fetch2_st,
		CU_0a_st,
		CU_0b_st,
		CU_1a_st,
		CU_1b_st,
		CU_2a_st,
		CU_2b_st,
		CU_3a_st,
		CU_3b_st,
		CU_4a_st,
		CU_4b_st,
		CU_5a_st,
		CU_5b_st,
		CU_6a_st,
		CU_6b_st,
		CU_7a_st,
		CU_7b_st,
		CU_8a_st,
		CU_8b_st,
		CU_9a_st,
		CU_9b_st,
		CU_10a_st,
		CU_10b_st,
		CU_11a_st,
		CU_11b_st,
		CU_12a_st,
		CU_12b_st,
		CU_13a_st,
		CU_13b_st,
		CU_idle1_st,
		CU_idle2_st
	);

	type tv_micro_codes is array (0 to 13) of std_logic_vector(41 downto 0);
	--Instruction Allocation--
	constant c_fetch      : tv_micro_codes := ("000000000000000000000100000000000100000000", "000000000000000000000001010000000000000000", "000000000000000000000000000000001000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) MI CO   (1) RO II       (2) CE
	constant c_LDA        : tv_micro_codes := ("000000000000000000000100100000000000000000", "000000000000000000000001001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) MI IO   (1) RO AI       (2) None					000001  LDA
	constant c_ADD        : tv_micro_codes := ("000000000000000000000100100000000000000000", "000000000000000000000001000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) MI IO   (1) RO BI       (2) AI EO FI				000010  ADD
	constant c_SUB        : tv_micro_codes := ("000000000000000000000100100000000000000000", "000000000000000000000001000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) MI IO   (1) RO BI       (2) AI EO SU FI			000011  SUB
	constant c_STA        : tv_micro_codes := ("000000000000000000000100100000000000000000", "000000000000000000000010000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) MI IO   (1) AO RI       (2) None					000100  STA
	constant c_LDI        : tv_micro_codes := ("000000000000000000000000101000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO AI   (1) None        (2) None					000101  LDI
	constant c_JMP        : tv_micro_codes := ("000000000000000000000000100000000010000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO CJ   (1) None        (2) None					000110  JMP / 00111 JMC / 01000 JMZ
	constant c_MOV_R0A    : tv_micro_codes := ("000000000000000000000000100000000000010000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R0AI (1) None        (2) None 					001001  MOV R0A
	constant c_MOV_R0B    : tv_micro_codes := ("000000000000000000000000100000000000001000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R0BI (1) None        (2) None					001010  MOV R0B
	constant c_MOV_R0     : tv_micro_codes := ("000000000000000000000000100000000000100000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R0I  (1) None        (2) None               001011  MOV R0
	constant c_MOV_A_R0A  : tv_micro_codes := ("000000000000000000000000001000000000000010", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R0AO (1) None        (2) None               001100  MOV A R0A
	constant c_MOV_A_R0B  : tv_micro_codes := ("000000000000000000000000001000000000000001", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R0BO (1) None        (2) None					001101  MOV A R0B
	constant c_OUT        : tv_micro_codes := ("000000000000000000000000000100010000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AO OI   (1) None        (2) None					001110  OUT
	constant c_HLT        : tv_micro_codes := ("000000000000000000001000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) HLT     (1) None        (2) None					001111  HLT
	constant c_MOV_A_R0   : tv_micro_codes := ("000000000000000000000000001000000000000100", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R0O  (1) None        (2) None					010000  MOV A R0
	constant c_MOV_R0_A   : tv_micro_codes := ("000000000000000000000000000100000000100000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AO R0I  (1) None        (2) None					010001  MOV R0 A
	constant c_MOV_R1A    : tv_micro_codes := ("000000000000000100000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R1AI (1) None        (2) None               010010  MOV R1A
	constant c_MOV_R1B    : tv_micro_codes := ("000000000000000010000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R1BI (1) None        (2) None               010011  MOV R1B
	constant c_MOV_R1     : tv_micro_codes := ("000000000000001000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R1I  (1) None        (2) None               010100  MOV R1
	constant c_MOV_A_R1A  : tv_micro_codes := ("000000000000000000100000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R1AO (1) None        (2) None               010101  MOV A R1A
	constant c_MOV_A_R1B  : tv_micro_codes := ("000000000000000000010000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R1BO (1) None        (2) None               010110  MOV A R1B
	constant c_MOV_A_R1   : tv_micro_codes := ("000000000000000001000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R1O  (1) None        (2) None               010111  MOV A R1
	constant c_MOV_R1_A   : tv_micro_codes := ("000000000000001000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AO R1I  (1) None        (2) None               011000  MOV R1 A
	constant c_MOV_R2A    : tv_micro_codes := ("000000000100000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R2AI (1) None        (2) None               011001  MOV R2A
	constant c_MOV_R2B    : tv_micro_codes := ("000000000010000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R2BI (1) None        (2) None               011010  MOV R2B
	constant c_MOV_R2     : tv_micro_codes := ("000000001000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO R2I  (1) None        (2) None               011011  MOV R2
	constant c_MOV_A_R2A  : tv_micro_codes := ("000000000000100000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R2AO (1) None        (2) None               011100  MOV A R2A
	constant c_MOV_A_R2B  : tv_micro_codes := ("000000000000010000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R2BO (1) None        (2) None               011101  MOV A R2B
	constant c_MOV_A_R2   : tv_micro_codes := ("000000000001000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AI R2O  (1) None        (2) None               011110  MOV A R2
	constant c_MOV_R2_A   : tv_micro_codes := ("000000001000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) AO R2I  (1) None        (2) None               011111  MOV R2 A
	constant c_ADD_R0A    : tv_micro_codes := ("000000000000000000000000000000100000000010", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R0AO BI (1) AI EO FI    (2) None					100000  ADD R0A
	constant c_ADD_R0B    : tv_micro_codes := ("000000000000000000000000000000100000000001", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R0BO BI (1) AI EO FI    (2) None					100001  ADD R0B
	constant c_ADD_R0     : tv_micro_codes := ("000000000000000000000000000000100000000100", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R0O BI  (1) AI EO FI    (2) None					100010  ADD R0
	constant c_SUB_R0A    : tv_micro_codes := ("000000000000000000000000000000100000000010", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R0AO BI (1) AI EO SU FI (2) None					100011  SUB R0A
	constant c_SUB_R0B    : tv_micro_codes := ("000000000000000000000000000000100000000001", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R0BO BI (1) AI EO SU FI (2) None					100100  SUB R0B
	constant c_SUB_R0     : tv_micro_codes := ("000000000000000000000000000000100000000100", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R0O BI  (1) AI EO SU FI (2) None					100101  SUB R0
	constant c_ADD_R1A    : tv_micro_codes := ("000000000000000000100000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R1AO BI (1) AI EO FI    (2) None               100110  ADD R1A
	constant c_ADD_R1B    : tv_micro_codes := ("000000000000000000010000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R1BO BI (1) AI EO FI    (2) None               100111  ADD R1B
	constant c_ADD_R1     : tv_micro_codes := ("000000000000000001000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R1O BI  (1) AI EO FI    (2) None               101000  ADD R1
	constant c_SUB_R1A    : tv_micro_codes := ("000000000000000000100000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R1AO BI (1) AI EO SU FI (2) None               101001  SUB R1A
	constant c_SUB_R1B    : tv_micro_codes := ("000000000000000000010000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R1BO BI (1) AI EO SU FI (2) None               101010  SUB R1B
	constant c_SUB_R1     : tv_micro_codes := ("000000000000000001000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R1O BI  (1) AI EO SU FI (2) None               101011  SUB R1
	constant c_ADD_R2A    : tv_micro_codes := ("000000000000100000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R2AO BI (1) AI EO FI    (2) None               101100  ADD R2A
	constant c_ADD_R2B    : tv_micro_codes := ("000000000000010000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R2BO BI (1) AI EO FI    (2) None               101101  ADD R2B
	constant c_ADD_R2     : tv_micro_codes := ("000000000001000000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R2O BI  (1) AI EO FI    (2) None               101110  ADD R2
	constant c_SUB_R2A    : tv_micro_codes := ("000000000000100000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R2AO BI (1) AI EO SU FI (2) None               101111  SUB R2A
	constant c_SUB_R2B    : tv_micro_codes := ("000000000000010000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R2BO BI (1) AI EO SU FI (2) None               110000  SUB R2B
	constant c_SUB_R2     : tv_micro_codes := ("000000000001000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) R2O BI  (1) AI EO SU FI (2) None               110001  SUB R2
	constant c_SET_P0x    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000010000000000000000001000000000000000", "000001000000000000000000001000000000000000", "000000100000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO BI   (1) P0O AI      (2) P0BO AI (3) AO P0I 110010 SET P0.x
	constant c_CLR_P0x    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000010000000000000000001000000000000000", "000011000000000000000000001000000000000000", "000000100000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) IO BI   (1) P0O AI      (2) P0BO CLR AI (3) AO P0I 110011 CLR P0.x
	constant c_MOV_A_P0   : tv_micro_codes := ("000000010000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) P0O AI  (1) None        (2) None        (3) None   110100 MOV A P0
	constant c_MOV_P0_A   : tv_micro_codes := ("000000100000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) P0I AO  (1) None        (2) None        (3) None   110101 MOV P0 A
	constant c_MOV_P0     : tv_micro_codes := ("000000100000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) P0I IO  (1) None        (2) None        (3) None   110110 MOV P0
	constant c_J_TF0      : tv_micro_codes := ("000000000000000000000000100000000011000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) TR0E IO CJ  FI (1) None   (2) None			 (3) None   110111  JB TF0 / 111000 JNB TF0
	constant c_S_C_T0E    : tv_micro_codes := ("100000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) T0E 	  (1) None			(2) None			 (3) None   111001 SET T0E / 111010 CLR T0
	constant c_MOV_TH0    : tv_micro_codes := ("001000000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) TH0I IO (1) None			(2) None			 (3) None   111100 MOV TH0
	constant c_MOV_TL0    : tv_micro_codes := ("000100000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) TL0I IO (1) None			(2) None        (3) None   111101 MOV TL0
	constant c_MOV_CS0    : tv_micro_codes := ("010000000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000"); -- (0) CS0I IO (1) None        (2) None        (3) None   111110 MOV CS0
	constant c_INC_R0A    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000010", "000000000000000000000000001010000001000000", "000000000000000000000000000100000000010000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R0B    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000001", "000000000000000000000000001010000001000000", "000000000000000000000000000100000000001000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R0     : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000100", "000000000000000000000000001010000001000000", "000000000000000000000000000100000000100000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R1A    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000100000001000000000000000", "000000000000000000000000001010000001000000", "000000000000000100000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R1B    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000010000001000000000000000", "000000000000000000000000001010000001000000", "000000000000000010000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R1     : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000001000000001000000000000000", "000000000000000000000000001010000001000000", "000000000000001000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R2A    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000100000000000001000000000000000", "000000000000000000000000001010000001000000", "000000000100000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R2B    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000010000000000001000000000000000", "000000000000000000000000001010000001000000", "000000000010000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R2     : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000001000000000000001000000000000000", "000000000000000000000000001010000001000000", "000000001000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R0A    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000010", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000010000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R0B    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000001", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000001000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R0     : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000100", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000100000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R1A    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000100000001000000000000000", "000000000000000000000000001011000001000000", "000000000000000100000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R1B    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000010000001000000000000000", "000000000000000000000000001011000001000000", "000000000000000010000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R1     : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000001000000001000000000000000", "000000000000000000000000001011000001000000", "000000000000001000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R2A    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000100000000000001000000000000000", "000000000000000000000000001011000001000000", "000000000100000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R2B    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000010000000000001000000000000000", "000000000000000000000000001011000001000000", "000000000010000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R2     : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000001000000000000001000000000000000", "000000000000000000000000001011000001000000", "000000001000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R0A   : tv_micro_codes := ("000000000000000000000000001000000000000010", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000010000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R0B   : tv_micro_codes := ("000000000000000000000000001000000000000001", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000001000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R0    : tv_micro_codes := ("000000000000000000000000001000000000000100", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000100000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R1A   : tv_micro_codes := ("000000000000000000100000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000100000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R1B   : tv_micro_codes := ("000000000000000000010000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000010000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R1    : tv_micro_codes := ("000000000000000001000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000001000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R2A   : tv_micro_codes := ("000000000000100000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000100000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R2B   : tv_micro_codes := ("000000000000010000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000010000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R2    : tv_micro_codes := ("000000000001000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000001000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_CALL       : tv_micro_codes := ("000000000000000000000000000000000100000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_RET        : tv_micro_codes := ("000000000000000000000000000000000010000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_PUSH_R0    : tv_micro_codes := ("000000000000000000000000000000000000000100", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_POP_R0     : tv_micro_codes := ("000000000000000000000000000000000000100000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_PUSH_R1    : tv_micro_codes := ("000000000000000001000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_POP_R1     : tv_micro_codes := ("000000000000001000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_PUSH_R2    : tv_micro_codes := ("000000000001000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_POP_R2     : tv_micro_codes := ("000000001000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DIR_P0     : tv_micro_codes := ("000000000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_JB_NB_P0_X : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000100000100000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000011000001000000", "000000000000000000000100000000000100000000", "000000000000000000000001000000000010000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_R3     : tv_micro_codes := ("000000000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_R3   : tv_micro_codes := ("000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_R3_A   : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_DM     : tv_micro_codes := ("000000000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_DM   : tv_micro_codes := ("000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_DM_A   : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MUL_R0     : tv_micro_codes := ("000000000000000000000000000000000000000000", "000000000000000000000000001000000000000100", "000000000000000000000000000000100000000000", "000000000000000000000000000011000001000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000000000000", "000000000000000000000000001000000000000100", "000000000000000000000000000000100000000000", "000000000000000000000000000011000001100000", "000000000000000000000000001000000000000000");
	constant c_DIV_R0     : tv_micro_codes := ("000000000000000000000000000000100000000100", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000001010000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MUL_R1     : tv_micro_codes := ("000000000000000000000000000000000000000000", "000000000000000001000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000011000001000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000000000000", "000000000000000001000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000001000000000000011000001000000", "000000000000000000000000001000000000000000");
	constant c_DIV_R1     : tv_micro_codes := ("000000000000000001000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000001010000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MUL_R2     : tv_micro_codes := ("000000000000000000000000000000000000000000", "000000000001000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000011000001000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000000000000", "000000000001000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000001000000000000000000011000001000000", "000000000000000000000000001000000000000000");
	constant c_DIV_R2     : tv_micro_codes := ("000000000001000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000001010000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_AND_R0     : tv_micro_codes := ("000000000000000000000000000000100000000100", "000011000000000000000000000000100000000000", "000011000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_AND_R1     : tv_micro_codes := ("000000000000000001000000000000100000000000", "000011000000000000000000000000100000000000", "000011000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_AND_R2     : tv_micro_codes := ("000000000001000000000000000000100000000000", "000011000000000000000000000000100000000000", "000011000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_AND_R3     : tv_micro_codes := ("000000000000000000000000000000100000000000", "000011000000000000000000000000100000000000", "000011000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_OR_R0      : tv_micro_codes := ("000000000000000000000000000000100000000100", "000001000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_OR_R1      : tv_micro_codes := ("000000000000000001000000000000100000000000", "000001000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_OR_R2      : tv_micro_codes := ("000000000001000000000000000000100000000000", "000001000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_OR_R3      : tv_micro_codes := ("000000000000000000000000000000100000000000", "000001000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_CPL_A      : tv_micro_codes := ("000000000000000000000000000100100000000000", "000000000000000000000000101000000000000000", "000011000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_XR0  : tv_micro_codes := ("000000000000000000000100000000000000000100", "000000000000000000000001001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_XR1  : tv_micro_codes := ("000000000000000001000100000000000000000000", "000000000000000000000001001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_XR2  : tv_micro_codes := ("000000000001000000000100000000000000000000", "000000000000000000000001001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_XR3  : tv_micro_codes := ("000000000000000000000100000000000000000000", "000000000000000000000001001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_XR0_A  : tv_micro_codes := ("000000000000000000000100000000000000000100", "000000000000000000000010000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_XR1_A  : tv_micro_codes := ("000000000000000001000100000000000000000000", "000000000000000000000010000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_XR2_A  : tv_micro_codes := ("000000000001000000000100000000000000000000", "000000000000000000000010000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_XR3_A  : tv_micro_codes := ("000000000000000000000100000000000000000000", "000000000000000000000010000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_INC_R3     : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DEC_R3     : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DJNZ_R3    : tv_micro_codes := ("000000000000000000000000001000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000010000001000000", "000000000000000000000000100000000010000000", "000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_ADD_R3     : tv_micro_codes := ("000000000000000000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SUB_R3     : tv_micro_codes := ("000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_P0x_C  : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000101000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000011100001000000", "000000010000000000000000001000000000000000", "000000000000000000000000100000100000000000", "000001100000000000000000000000000000000000", "000011100000000000000000000000000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_C_P0x  : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000100000000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000100000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_RDA_P0     : tv_micro_codes := ("000000000000000000000000100000000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_ADDI       : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SUBI       : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_DIR_P1     : tv_micro_codes := ("000000000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_P1     : tv_micro_codes := ("000000000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_P1_A   : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_P1   : tv_micro_codes := ("000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SET_P1x    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000000", "000001000000000000000000001000000000000000", "000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_CLR_P1x    : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001000000000000000", "000011000000000000000000001000000000000000", "000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_P1x_C  : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000101000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000100000000000", "000000000000000000000000000011100001000000", "000000000000000000000000001000000000000000", "000000000000000000000000100000100000000000", "000001000000000000000000000000000000000000", "000011000000000000000000000000000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_C_P1x  : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000100000000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000100000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_RDA_P1     : tv_micro_codes := ("000000000000000000000000100000000000000000", "000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_CMPI       : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000000011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_CMP        : tv_micro_codes := ("000000000000000000000100100000000000000000", "000000000000000000000001000000100000000000", "000000000000000000000000000011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_TH0_A  : tv_micro_codes := ("001000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_TL0_A  : tv_micro_codes := ("000100000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_CS0_A  : tv_micro_codes := ("010000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_TC0L : tv_micro_codes := ("000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_TC0H : tv_micro_codes := ("000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SET_TCR0E  : tv_micro_codes := ("000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_JB_NB_T0V  : tv_micro_codes := ("000000000000000000000000100000000010000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_PC_A   : tv_micro_codes := ("000000000000000000000000000100000010000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_PC   : tv_micro_codes := ("000000000000000000000000001000000100000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_LR     : tv_micro_codes := ("000000000000000000000000100000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_LR_A   : tv_micro_codes := ("000000000000000000000000000100000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_A_LR   : tv_micro_codes := ("000000000000000000000000001000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_PC_LR  : tv_micro_codes := ("000000000000000000000000000000000010000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_MOV_LR_PC  : tv_micro_codes := ("000000000000000000000000000000000100000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SUBB_R0    : tv_micro_codes := ("000000000000000000000000000000100000000100", "000000000000000000000000001011000001000000", "000000000000000000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SUBB_R1    : tv_micro_codes := ("000000000000000001000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SUBB_R2    : tv_micro_codes := ("000000000001000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SUBB_R3    : tv_micro_codes := ("000000000000000000000000000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SUBIB      : tv_micro_codes := ("000000000000000000000000100000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	constant c_SUBB       : tv_micro_codes := ("000000000000000000000100100000000000000000", "000000000000000000000001000000100000000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000100000000000", "000000000000000000000000001010000001000000", "000000000000000000000000001011000001000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000");
	

	constant cv_IC_NOP		  : std_logic_vector := X"00";
	constant cv_IC_LDA        : std_logic_vector := X"01";
	constant cv_IC_ADD        : std_logic_vector := X"02";
	constant cv_IC_SUB        : std_logic_vector := X"03";
	constant cv_IC_STA        : std_logic_vector := X"04";
	constant cv_IC_LDI        : std_logic_vector := X"05";
	constant cv_IC_JMP        : std_logic_vector := X"06";
	constant cv_IC_JMC        : std_logic_vector := X"07";
	constant cv_IC_JMZ        : std_logic_vector := X"08";
	constant cv_IC_MOV_R0A    : std_logic_vector := X"09";
	constant cv_IC_MOV_R0B    : std_logic_vector := X"0a";
	constant cv_IC_MOV_R0     : std_logic_vector := X"0b";
	constant cv_IC_MOV_A_R0A  : std_logic_vector := X"0c";
	constant cv_IC_MOV_A_R0B  : std_logic_vector := X"0d";
	constant cv_IC_OUT        : std_logic_vector := X"0e";
	constant cv_IC_HLT        : std_logic_vector := X"0f";
	constant cv_IC_MOV_A_R0   : std_logic_vector := X"10";
	constant cv_IC_MOV_R0_A   : std_logic_vector := X"11";
	constant cv_IC_MOV_R1A    : std_logic_vector := X"12";
	constant cv_IC_MOV_R1B    : std_logic_vector := X"13";
	constant cv_IC_MOV_R1     : std_logic_vector := X"14";
	constant cv_IC_MOV_A_R1A  : std_logic_vector := X"15";
	constant cv_IC_MOV_A_R1B  : std_logic_vector := X"16";
	constant cv_IC_MOV_A_R1   : std_logic_vector := X"17";
	constant cv_IC_MOV_R1_A   : std_logic_vector := X"18";
	constant cv_IC_MOV_R2A    : std_logic_vector := X"19";
	constant cv_IC_MOV_R2B    : std_logic_vector := X"1a";
	constant cv_IC_MOV_R2     : std_logic_vector := X"1b";
	constant cv_IC_MOV_A_R2A  : std_logic_vector := X"1c";
	constant cv_IC_MOV_A_R2B  : std_logic_vector := X"1d";
	constant cv_IC_MOV_A_R2   : std_logic_vector := X"1e";
	constant cv_IC_MOV_R2_A   : std_logic_vector := X"1f";
	constant cv_IC_ADD_R0A    : std_logic_vector := X"20";
	constant cv_IC_ADD_R0B    : std_logic_vector := X"21";
	constant cv_IC_ADD_R0     : std_logic_vector := X"22";
	constant cv_IC_SUB_R0A    : std_logic_vector := X"23";
	constant cv_IC_SUB_R0B    : std_logic_vector := X"24";
	constant cv_IC_SUB_R0     : std_logic_vector := X"25";
	constant cv_IC_ADD_R1A    : std_logic_vector := X"26";
	constant cv_IC_ADD_R1B    : std_logic_vector := X"27";
	constant cv_IC_ADD_R1     : std_logic_vector := X"28";
	constant cv_IC_SUB_R1A    : std_logic_vector := X"29";
	constant cv_IC_SUB_R1B    : std_logic_vector := X"2a";
	constant cv_IC_SUB_R1     : std_logic_vector := X"2b";
	constant cv_IC_ADD_R2A    : std_logic_vector := X"2c";
	constant cv_IC_ADD_R2B    : std_logic_vector := X"2d";
	constant cv_IC_ADD_R2     : std_logic_vector := X"2e";
	constant cv_IC_SUB_R2A    : std_logic_vector := X"2f";
	constant cv_IC_SUB_R2B    : std_logic_vector := X"30";
	constant cv_IC_SUB_R2     : std_logic_vector := X"31";
	constant cv_IC_SET_P0X    : std_logic_vector := X"32";
	constant cv_IC_CLR_P0X    : std_logic_vector := X"33";
	constant cv_IC_MOV_A_P0   : std_logic_vector := X"34";
	constant cv_IC_MOV_P0_A   : std_logic_vector := X"35";
	constant cv_IC_MOV_P0     : std_logic_vector := X"36";
	constant cv_IC_JB_TF0     : std_logic_vector := X"37";
	constant cv_IC_JNB_TF0    : std_logic_vector := X"38";
	constant cv_IC_SET_T0E    : std_logic_vector := X"39";
	constant cv_IC_CLR_T0     : std_logic_vector := X"3a";
	constant cv_IC_SET_TR0    : std_logic_vector := X"3b";
	constant cv_IC_MOV_TH0    : std_logic_vector := X"3c";
	constant cv_IC_MOV_TL0    : std_logic_vector := X"3d";
	constant cv_IC_MOV_CS0    : std_logic_vector := X"3e";
	constant cv_IC_INC_R0A    : std_logic_vector := X"3f";
	constant cv_IC_INC_R0B    : std_logic_vector := X"40";
	constant cv_IC_INC_R0     : std_logic_vector := X"41";
	constant cv_IC_INC_R1A    : std_logic_vector := X"42";
	constant cv_IC_INC_R1B    : std_logic_vector := X"43";
	constant cv_IC_INC_R1     : std_logic_vector := X"44";
	constant cv_IC_INC_R2A    : std_logic_vector := X"45";
	constant cv_IC_INC_R2B    : std_logic_vector := X"46";
	constant cv_IC_INC_R2     : std_logic_vector := X"47";
	constant cv_IC_DEC_R0A    : std_logic_vector := X"48";
	constant cv_IC_DEC_R0B    : std_logic_vector := X"49";
	constant cv_IC_DEC_R0     : std_logic_vector := X"4a";
	constant cv_IC_DEC_R1A    : std_logic_vector := X"4b";
	constant cv_IC_DEC_R1B    : std_logic_vector := X"4c";
	constant cv_IC_DEC_R1     : std_logic_vector := X"4d";
	constant cv_IC_DEC_R2A    : std_logic_vector := X"4e";
	constant cv_IC_DEC_R2B    : std_logic_vector := X"4f";
	constant cv_IC_DEC_R2     : std_logic_vector := X"50";
	constant cv_IC_DJNZ_R0A   : std_logic_vector := X"51";
	constant cv_IC_DJNZ_R0B   : std_logic_vector := X"52";
	constant cv_IC_DJNZ_R0    : std_logic_vector := X"53";
	constant cv_IC_DJNZ_R1A   : std_logic_vector := X"54";
	constant cv_IC_DJNZ_R1B   : std_logic_vector := X"55";
	constant cv_IC_DJNZ_R1    : std_logic_vector := X"56";
	constant cv_IC_DJNZ_R2A   : std_logic_vector := X"57";
	constant cv_IC_DJNZ_R2B   : std_logic_vector := X"58";
	constant cv_IC_DJNZ_R2    : std_logic_vector := X"59";
	constant cv_IC_CALL       : std_logic_vector := X"5a";
	constant cv_IC_RET        : std_logic_vector := X"5b";
	constant cv_IC_PUSH_R0    : std_logic_vector := X"5c";
	constant cv_IC_POP_R0     : std_logic_vector := X"5d";
	constant cv_IC_PUSH_R1    : std_logic_vector := X"5e";
	constant cv_IC_POP_R1     : std_logic_vector := X"5f";
	constant cv_IC_PUSH_R2    : std_logic_vector := X"60";
	constant cv_IC_POP_R2     : std_logic_vector := X"61";
	constant cv_IC_DDRP0      : std_logic_vector := X"62";
	constant cv_IC_JB_P0x     : std_logic_vector := X"63";
	constant cv_IC_JNB_P0x    : std_logic_vector := X"64";
	constant cv_IC_JB_P1x     : std_logic_vector := X"65";
	constant cv_IC_JNB_P1x    : std_logic_vector := X"66";
	constant cv_IC_MOV_R3     : std_logic_vector := X"73";
	constant cv_IC_MOV_A_R3   : std_logic_vector := X"74";
	constant cv_IC_MOV_R3_A   : std_logic_vector := X"75";
	constant cv_IC_MOV_DM     : std_logic_vector := X"76";
	constant cv_IC_MOV_A_DM   : std_logic_vector := X"77";
	constant cv_IC_MOV_DM_A   : std_logic_vector := X"78";
	constant cv_IC_MUL_R0     : std_logic_vector := X"79";
	constant cv_IC_DIV_R0     : std_logic_vector := X"7a";
	constant cv_IC_MUL_R1     : std_logic_vector := X"7b";
	constant cv_IC_DIV_R1     : std_logic_vector := X"7c";
	constant cv_IC_MUL_R2     : std_logic_vector := X"7d";
	constant cv_IC_DIV_R2     : std_logic_vector := X"7e";
	constant cv_IC_PUSH_DM    : std_logic_vector := X"7f";
	constant cv_IC_POP_DM     : std_logic_vector := X"80";
	constant cv_IC_PUSH_R3    : std_logic_vector := X"81";
	constant cv_IC_POP_R3     : std_logic_vector := X"82";
	constant cv_IC_AND_R0     : std_logic_vector := X"83";
	constant cv_IC_AND_R1     : std_logic_vector := X"84";
	constant cv_IC_AND_R2     : std_logic_vector := X"85";
	constant cv_IC_AND_R3     : std_logic_vector := X"86";
	constant cv_IC_OR_R0      : std_logic_vector := X"87";
	constant cv_IC_OR_R1      : std_logic_vector := X"88";
	constant cv_IC_OR_R2      : std_logic_vector := X"89";
	constant cv_IC_OR_R3      : std_logic_vector := X"8a";
	constant cv_IC_CPL_A      : std_logic_vector := X"8b";
	constant cv_IC_MOV_A_atR0 : std_logic_vector := X"8c";
	constant cv_IC_MOV_A_atR1 : std_logic_vector := X"8d";
	constant cv_IC_MOV_A_atR2 : std_logic_vector := X"8e";
	constant cv_IC_MOV_A_atR3 : std_logic_vector := X"8f";
	constant cv_IC_MOV_atR0_A : std_logic_vector := X"90";
	constant cv_IC_MOV_atR1_A : std_logic_vector := X"91";
	constant cv_IC_MOV_atR2_A : std_logic_vector := X"92";
	constant cv_IC_MOV_atR3_A : std_logic_vector := X"93";
	constant cv_IC_INC_R3     : std_logic_vector := X"94";
	constant cv_IC_DEC_R3     : std_logic_vector := X"95";
	constant cv_IC_DJNZ_R3    : std_logic_vector := X"96";
	constant cv_IC_ADD_R3     : std_logic_vector := X"97";
	constant cv_IC_SUB_R3     : std_logic_vector := X"98";
	constant cv_IC_MOV_P0X_C  : std_logic_vector := X"99";
	constant cv_IC_MOV_C_P0X  : std_logic_vector := X"9a";
	constant cv_IC_RDA_P0     : std_logic_vector := X"9b";
	constant cv_IC_MOV_A_C    : std_logic_vector := X"9c";
	constant cv_IC_MOV_C_A    : std_logic_vector := X"9d";
	constant cv_IC_MOV_C      : std_logic_vector := X"9e";
	constant cv_IC_RRC        : std_logic_vector := X"9f";
	constant cv_IC_RLC        : std_logic_vector := X"a0";
	constant cv_IC_PUSH_A     : std_logic_vector := X"a1";
	constant cv_IC_POP_A      : std_logic_vector := X"a2";
	constant cv_IC_ADDI       : std_logic_vector := X"a3";
	constant cv_IC_SUBI       : std_logic_vector := X"a4";
	constant cv_IC_DDRP1      : std_logic_vector := X"b5";
	constant cv_IC_MOV_P1     : std_logic_vector := X"b6";
	constant cv_IC_MOV_P1_A   : std_logic_vector := X"b7";
	constant cv_IC_MOV_A_P1   : std_logic_vector := X"b8";
	constant cv_IC_SET_P1X    : std_logic_vector := X"b9";
	constant cv_IC_CLR_P1X    : std_logic_vector := X"ba";
	constant cv_IC_MOV_P1X_C  : std_logic_vector := X"bb";
	constant cv_IC_MOV_C_P1X  : std_logic_vector := X"bc";
	constant cv_IC_RDA_P1     : std_logic_vector := X"bd";
	constant cv_IC_CMPI       : std_logic_vector := X"be";
	constant cv_IC_CMP        : std_logic_vector := X"bf";
	constant cv_IC_MOV_A_TH0  : std_logic_vector := X"c0";
	constant cv_IC_MOV_A_TL0  : std_logic_vector := X"c1";
	constant cv_IC_MOV_CS0_A  : std_logic_vector := X"c2";
	constant cv_IC_ADDC_R0    : std_logic_vector := X"c3";
	constant cv_IC_ADDC_R1    : std_logic_vector := X"c4";
	constant cv_IC_ADDC_R2    : std_logic_vector := X"c5";
	constant cv_IC_ADDC_R3    : std_logic_vector := X"c6";
	constant cv_IC_ADDIC      : std_logic_vector := X"c7";
	constant cv_IC_ADDC       : std_logic_vector := X"c8";
	constant cv_IC_MOV_A_TC0L : std_logic_vector := X"c9";
	constant cv_IC_MOV_A_TC0H : std_logic_vector := X"ca";
	constant cv_IC_SET_TCR0E  : std_logic_vector := X"cb";
	constant cv_IC_JB_T0V     : std_logic_vector := X"cc";
	constant cv_IC_JNB_T0V    : std_logic_vector := X"cd";
	constant cv_IC_SET_TC0L   : std_logic_vector := X"ce";
	constant cv_IC_MOV_PC_A   : std_logic_vector := X"cf";
	constant cv_IC_MOV_A_PC   : std_logic_vector := X"d0";
	constant cv_IC_MOV_LR     : std_logic_vector := X"d1";
	constant cv_IC_MOV_LR_A   : std_logic_vector := X"d2";
	constant cv_IC_MOV_A_LR   : std_logic_vector := X"d3";
	constant cv_IC_MOV_PC_LR  : std_logic_vector := X"d4";
	constant cv_IC_MOV_LR_PC  : std_logic_vector := X"d5";
	constant cv_IC_SUBB_R0    : std_logic_vector := X"d6";
	constant cv_IC_SUBB_R1    : std_logic_vector := X"d7";
	constant cv_IC_SUBB_R2    : std_logic_vector := X"d8";
	constant cv_IC_SUBB_R3    : std_logic_vector := X"d9";
	constant cv_IC_SUBIB      : std_logic_vector := X"da";
	constant cv_IC_SUBB       : std_logic_vector := X"db";
	

	constant ci_max_control_L : integer := 69;

end control_fsm_p;
